/**
 * @Author: Qiao Zhang
 * @Date: 2025-12-18 22:21:47
 * @LastEditTime: 2026-01-01 20:56:27
 * @LastEditors: Qiao Zhang
 * @Description: Some important definitions which will be shared in different files
 * @FilePath: /cnn/hardware/rtl/include/definitions.sv
 */

`ifndef DEFINITIONS
    `define DEFINITIONS
    `timescale 1ns/1ps
    package definitions;

        // ==========================================================
        //  1.  Global Hardware Specs (Synthesized Constants)
        // ==========================================================
        parameter int INT_WIDTH         = 8;

            // Max supported Kernel Size (e.g. 7x7), determines Pointer Pool size
        parameter int MAX_K_R           = 7;

            // Line Buffer Depth: Supports full HD width
        parameter int MAX_LINE_W        = 1920;

            /*
                The Physical Width of the Systolic Array / ARR
                This is the "Modulo" basis for Circular Buffering.
                Even if Image is 1920 wide, we map it to these 64 columns.
            */
        parameter int MAX_TILE_W        = 64;

        // ==========================================================
        // 2. Model Default Parameters (Can be overridden by Software Config)
        // ==========================================================

        parameter int K_CHANNELS        = 6;

            // A. Systolic Arrays IP
                // Mode 0: save area(just 1 adder for 1 pe --- blocking)
                // Mode 1: high performance(multi adder for 1 pe --- non-blocking, pipeline)
        parameter int MODE         = 0              ;

        parameter int MATRIX_A_ROW = K_CHANNELS     ;
        parameter int MATRIX_A_COL = 25             ;
        parameter int MATRIX_B_ROW = MATRIX_A_COL   ;
                // NOTE: Systolic Array Columns.
                // If MAX_TILE_W (64) > MATRIX_B_COL (16), the Wrapper manages the mapping.
        parameter int MATRIX_B_COL = 64             ;
        parameter int DATA_WIDTH   = INT_WIDTH      ;
        parameter int ACC_WIDTH    = 32             ;

            // B. column_fifo
        parameter int COLUMN_FIFO_DEPTH = 8         ;// Enough for 5x5 or 7x7

            // C. Input_buffer_bank
                // Instantiates enough FIFOs to hold a FULL HD Line
        parameter int IB_BANK_W         = MAX_LINE_W;

            // D. Active Row Register
        parameter int PTR_WIDTH         = 32;  // the pre-wave pointer width

            // E. Global Buffer
        parameter int SRAM_DEPTH        = 4096      ;// 4kB
        parameter int SRAM_ADDR_W       = $clog2(SRAM_DEPTH);

    endpackage
    import definitions::*;
`endif
